BZh91AY&SY%?�q l`߀py����������`K�|�AQ��Q�T��HR�s�}��Ǣ+jJ�������ݲJ�����L��u�(�2R��(��7Mh������J�n����i���� �3���P�Q�\��YV��歛dؑި      ��Rm��T�(i�J�I�@ ���2 ɦ���"��z��F�  ���� �)IT��4hѠ      i"E$�2h      )JI�3H�S2��&M=#�d�# CM4$!  	��S��MOFS���4�h�M9��=U9s�� ��;�Sa *�����z�!U7Ɨ�{)Ok��je�)��J֓�U Z*���RI?�tA5�ȉ��H@��z�=��Oy]��G_g�����[ۣ}�O�gLL:at�qS4Q�Q���H�B3i��D"0�#6�����E�da��شQE5h����#�P�L�4�����i:�e3*����!�C��RE2I�(�"�F�RQ!F���T���"�>0�5h]*�1?Di�#��F��[�AtF#�!}�VPDY��!��*e�eN��C,�E�H��]2�d2���ߍ�;�����	:eԿ�B(��^��͖B!�%@��uB!:�+K����Qt���	j�M^ �U'��{�La�-֑e*����"ZY����~��E"��
�vE�0�"&L��}F��!6�FGЈa�>�Bd��U�hU�#DQ���"����d���!�+�#�u�|���L{�mi�du�|�/��͐�����2Ϟ�"*͡d�L�2B>W^D~�l����>�!�B�C�}"ԅe?�1S��)���g!�6������S�U~F�(���0�>��#���`qY}�Јa&Z���G�F8Ցg̊"@�B!򢊪��l9�~̼9�A�Xe�ƑJ���(��gC���/Qx-�7U��y�@e�p� �}�%URI����f���]г�"̒O�!���\m��׌��2�G��F:�1��^���_t�}��(����sX�k�F��}�&i�J�G��~����jƩ����%hU@�,�1�FD	�,�Ą����@�Y�lZ%����r��i@B"�g[�P?ge��ڰ�*�����$v܊����3���2���̼e^O��F�A��E�l�n��m@A�v���	�Fc9���*��{$����ʴb�DO#�h9|j��W5u��*8�\\O%��Xg'J��dp�W�w�a��,����:0׆���#R
�4��:��m ����_��N��P���-�S)�7����ئr�;r�&�-ڛ]�Ic͈(�j���Z�l�6(�s�p�7���.�f�^]ϳH��H�V��+�a��sEX'm��e5V���Wk�/7V+7w54���7Bƕ��睮�s֘qPN�
���/2� �Kdo���'�V,�"*��*���7�ŗe�O�.��v1Ian`�)V>Da�`���rԨ��a����Y ��@�B��![�IR8�3d�|�N��R��+�]�/�mR�>6�I��[�A�X�U�N��ԣVB�&�/��»x��N��В��=w���J��L;r�գ3yuS� ��fȽ"l�s�8l90�y۴�%��e؊�f���-��W��\��w���
���3g;/8�铛�6�A\m�w�-V6≤l�d	��N�e���}nesp���$�t�yb���4���b]ܷ�*##gT���%��Y�^J>�}Ec���nuPSb֕CӮ�5��'5�k�n��sv�����%a�{8Yaj�zݞ�{����Ujj��Hb����b/����Rʁ�a	ūҗwM뫿\2-�8R�.��f���wf�h�Y�E[F���!~�J��4���3.[�rU9WG�Q��h>���2�氭��0ĕ�{��>�u�l���[��Л��;0%�][R�@M^��G�*�۫4�kǺ	�cH�L=���6ƭ��J�{;�6Gy�m��8J�r�}z�ַ��xGky`{�Ye)\ҕafɧMAPUC3�H�2�!�$Ȅ��̵[��F(�e�e��i��n�+Wlį���w�خTӒ��]W'��o����J[�1a�h���
��`��Ҿ�7�8 ԫ�oEV�3y��q!͚%J�t������:��{�u'Yn�7�ӠMj�|z^�2f�p���I��QXkn8�X<+��a�1at�+�v�[��^Wp�"缄��TۓU����YYz�:|n�N�0�K\�w8��ٰK���0�`�K�m�zFwt�o����Or��n�#D/B��I��>$�D6�ȺJoy��D��0��]���ݏ�ZSz,�iu�&��,��`o7��'n:���z����G)dW��`cN"1":ݔ���9����pv���%S/9k��(�����i�!���Y�6In=�X9�[nI|�<���̓Q͂�
�e���T�m�C��c&��ӧN�
h��$4}L �dT
$M1���[Tj�Q0�>�D�^1��H$��@��0"Q)�*�)���Q �X۶�H�L�H>>�LST�EO�M�r�b�B��U��Q	FۻlI�	-Ў"���HUOP��4A"�I�R ̪�9 �� �
��"��q3��Pā�,��#J����m�1+4��WM���+���ԹN5L�����Y������f���b��/(Q�כX���f<論��Y���1���i���6�TC30��k\]heQUYY:�*�-u�r�b���""W�f3XSV���*����m�[O�Tԇ?�0��!m[��U
Ēh����.6�}{d���5�}Y���������������Z����>��}:�>P�}G��O��{�.>��_K2H��owvwwvwwrI%)$�$�$�����K)$�Z�I$�H$�I$�I$��RI$�'I$���"RI$�K�J��I$�'I$���$�����R�J�JI+I(I$�$�$�ĊI$���I$�	$�I �)$�JC0)$� �I$�	$�KQI$�ĝ$�V���IZJI*I)I%)$�$�$�����J�N�I,H�)$�P������|}#�f,fHH:�r���u�G�U�7�-�Q�{}�����4�em��G�?����$�W�Mg��d���bm\5	 ��~��36�EY$��,ѤRO9�n�`]㨈�A��l����F)Ҵ7U�=S�\w�i�wv-K�k֯��r�\�=����g�a9����"bB\� �d6L�. ���NF$���c�l��vc�Ma��{)��ٯD�u�K/MS(�U���C9�y}�i����ԇP{�Q�@��mM�O��Ύ�:�7��1.d��-�z��k�ʶ�7w�1E�p���]A�����}a*�Q�z�Urq��n��~a���Ò~�#����$����pӦ�����Z����B�tU)5IF�)x����f4�h�j�9$�3��(�H��1���g3��U�U1���ߤ��]���=f<��3�����R��d�Jא�B>��Q�7%��߽�f�h�Cs�T{��c�3Z�;m�~7J�$���&�R+=*r4����g�iq�4��@�vS8�a6�8�!W8{�k�Q$��Y�{n����׽�"w�����h���*+�1��L��zd�{ۋֳxr�.��˪$��jro�	��$r�I�2�4<,�x�W�
uh;Ef���gv�G*�n;*�ZU6�$��E9`�z�]�B�Z�o���Ч��.�:�Ir��>�R"�!���Y$��]�G
��7BY�6oV�=�8�דS�y�4���d�s���Up�$�ܫ:w$��v/(�b>=�V���l�]=��ۏ5U�h��Z�g3j1b!hhe���AHT6�w&�&���W�-u!ru�?x'┘T������$���ǫkA��!Z�n��o�`�%����Zg��+jMȣO����UD�ٶ��*�r��nVԱ�5K���X��H��2Q`�σX�L#�"4���l&!4���cV�������aYN�F�M۽������"����ΰJ��f]��7V�A#�u�`鷓x3aKj�o`K�1�5�X7�iqDQr[���h�N�|����|�������~�����)C�I$�J8H���q%�t�=��J�I$���;sBc�,�g<���ȁ����`ވ|x8�QJ&F��4U��ﲽ6�e��	�UB>���$�3�u� t�_=/­���l��TA�_�ʵ�>qS�4����.&	G/ޠ�Q@�k�(��A���Y&��8�M�O蝚�J�?i@�C�4M$��ۦ`��p#2��+����H=X���1�}�0&I$�6���D��޻�Q������$��8��������uw���%�dF���"ֽF���dߢ�4}D�O�z�۠	H� at`,��c�3k���PW�Wͦ}�fK<Õ���i�(R��ұ;�f�-%4t�D�p��74:,m��I%P�����8����9f��g<_U��t�ºw���[��3P�#8%w�X���<��D;�#P���#��G|�&S�ߺY%�� ��xɮ/�-%�@����xq�x��c*�+��.-�;�6��F�Z4�5�p�x�I���8}��̗�	�(|8[_X��D���q>�����0�\��@Z.m�6a���soP1����8� "�1��p�8����?;[<	�r&D ]#z��3Zž n0����G�>0�kTG��Q�4�����x�AÜ�3( �C�X)�!}�'����G��8a�w����ޢ��`xHTEb��ij#1[��b����u�h��
m�"|?=(��;K��y���Q\�����^H�ɼ�P5���G)��7�YqL�b۹6�<����=X��(v��]e�F�O�@�뤀����B����6\�M2��3I�����~�g��:U�g����bIbI�D�I+I:� �)ٚ�hu�b<�=��1���E���ˣ� �9a����1�
s��a��-�mZ�E�,�YWP~�^]�\v��0= Գq�>�H���ٌ�6��šy>�㙃�s����գ6�жt0��@7EK�hE0^��[�I 	9�(U?_}��Sd�hn�F����=uF&��ΈX|���$IW�!s> ��!��cf�5el̠�y��ǹ|G�t��讛~�fɋ皨p 34�p�r��8��z�������Pe�B��y����xq�z�}e[\�"�h���=�ԇ���|t�u�@��f8i�`#3�	~�������a�N���z�����ܷt��DZ��z�/Jˋ�F@�L��<��DV��{~�h��dP�f�q��n��U�Q3V��0F,(�B�	���_�A��:��y�i$4�,� ��p�9�V�a
|9ـ�E���4����(���c�4O�����vE����S\4�Z�/{��-�7��~Z�����}gq��/������{��z 'qJ=;���gީ"j�@s:\a��cP���K!����b`qe0���:h��$W�=��a�b�𚰁� �!`q]�"x37-�~w�S��C�&���2�V.9��8�(����L�̰�Dy��j���r�v�$] D�\�����7�Ȍ�#���h���U*����p�*UJ���`=�0&���|�!��f�S4ENE�P=L8����p�d�ΐ6�t3��^  v�h��(�֥E��D�e��T(�(��EH��[JDx	���5C�}*P��JHC�*�)���K��|�4�$KV����W2����d�͛�{˹c*�6���.�^�]��r�^Ԇ��5�'j\���@;tz]��ܝDL$�������V�u0�J�J"��UT\[������7���¨��#�̼�����>�=�h�Κ�$0�����FR���8f�(!��i���3K��RE� �T����R����Z�f�S���82x��q�$,@z.I�30ʃ)q����h��]`i'.�4v�ڤ7���7ƣ���Ծ�_��N�#���6{ĳ����B��������~�T&s���F���.�>1�7�f�� �u ���m���z�K�k�bf�T�G";�^��y7��A�qWU.g�.�	�tj���<��
��C�i/.:F�;�~���<d�<��=4�r`9�a�q{�,�5yY��8M���� 0(9$mڡ��>��\fz!�p������<�
#���/{©M(|��n$դ8�S��Ԏ�?�a�ԍG>��GmR�C)��.�
?a�	CA`�#�S����X�Ȳ��LA�Op>$+���h�n�c�fT��	ۋ�'���A
ψß��5�fA�U"Î�cq�6g�]�enE���E�<=M	A�!�vzM���u���zO� �&�IE5�{�4q�x���|.#
�dCUM����}�J��Df�*�7�>�p� @����������H����N ��Ꮬ_@��f��r�Q.�=�>�7��j9�\�}�I ��(z�ネ'��OW��qL@hWV��J*��_���M��;݅jk~�o۬�[�ok�G6"��5����\볕�>��>��Tѯ1@�i�ܥ��rt����
1&�����	d�E����e�A" M�BE���m=�ͤ�����T�Q"RIRIGѹv`r��O�#�H�����	s�k(O���J��/�j�p�>{#���3�3�J�\�<���꫖��Ⴄ9ó�0{���7�Ќ�_�=�r��"~���//�͸dK��˹+\I&H�2�>`�/K�	��8��1�f��BCzc�֛����z"�ަ���h	���;�'��"��, ���O�~�凘4�Ȑ�|D+���Ӿ����w��Tut��N�8�ۇ�v
�\����G��,���Z��r����g���?���\�F�`�p8�^�>�0ϊ�ir�"'{1z�<����n���{C'wh��q�������s���4����݈�qdWxs�C�� �:�C��/�������d���AQ67u��x0K�r�N��@�:����Bp���r��N�:(����|�R����D_�P�(j�J������Ga�06������5��b�E���
Κ��^ݥ�wt�l<����n���:���5�(Y�	z�o�K
<l�ar���aϢboM#��/aϹ=�K�,�[���Et�vI���W;��rq��.Q&#��(�?��HSel��(>�2@��z��0�#�ᅑ'H�$E�ϋ*v��C��ހ���5Q�|��WNp���i� �Dа��<�]��O�l]3� e�]	����7��f�ya�PEru��a}ݒ��'Ҫ߾J�4�{�L��!c݉���+R�D�AƵ
�d�IFZ�R�)	"QD�챬S�y�W��N�����oY�s�AT�!�`H�B�Ym�N�j�0O�>�&'��>;ۯ,:כ�7�ml{19�Ȕ�i۳�s���!h�Ėz�c�o�0�sGQ��j�s�<�٬V����.]��F>4Aбa����
s�\�<��6��w��c��P���Oon���k�s5��jR=�b�r4`�j�z�#:�ژ�}ɔ��\չ[c������
�{+�wݗU����~]ٽ<���T�R�Q
�JRJ"!RIJIG0����^�
���_��ϐ/6�$�����΃&�g���x�hzNw�:O��d���gHk|��G��;���N?�Լ9l� a ��-�]$����0��*O�`���vvj��Caas1s=��p��E�LC�/S���/�m����������\�s��h����E���~�kU #����-�8.�\�z�j<�c���Y[��l��0g36�U^���� {<�vs�)�i�Ͳ��r��m���.T�(Iw�����Ey����ǮzE��0�Fhf`*w����ٮ$�Ӕ8ƻ�N ��	$1�ѽ.]����^4	�a�
"HD�Ȃ>�q�b�|�qs�5�ia��1s^y"�(
	��+tsKטK4$�T����T�����<r���8r8y��LΜ��[�z�c	0��d��g#�?ǭ�[I�P��M�/>^�z q����yt�N]ށ81e�Lo���J���Q���$x�kz�����&1�,v(˔Q������ps����Zb�4��l74!�~��u �XJv��9�Y:ss˼���Q���NS�������ǚĔq}�U�L��P{��W���M5���s�=.�x�M%�F�o��l��L՚�5E��T���b���g%�Tb�Q|ҬR�"��4��{�4��S-�� �ʲ���[R#	�B����i���o�N˓2��v�Ǝ�/{%h�U�M��*&y3�
�z��e��`��6K���lޜ#�o���
[������/v"K��D.D2�R���d�h��JM=�n�	'wIZJN�$����Yh>�M&����4v�����Ѡ���wosP�����UwV��-�� (�5�͸��wG���6���3�������!�6�õf��`�qO&��:"A*�G���V�b�u!s0��VH�D.�9ۤ��f��73�T		ǽ�	%�W'G3�y�3?<��)�G�*v2}��)�æ��pX,�W�y�8ffܽS; �^����^���=�R�G�m:3�V����l������� a�n��l�`=M������!�'&]ܯD��4��o:G�1����%育����$)̥jG�K, ���yx��LS0`6��}�&�T)�6�%���D�0բ�������0�f�|Y������������5��Ӭ��5���n�*!�>f�È|lH�<`U����<4�j�P����1����3����h�"�ס�j6�YN���O��w5f���uq+�<���l��` 
���^����&cA���P�q�r�㞕[��.N]8�n���Jp�al^��y�t�ḫ�ܘ;
5����a�;�HԳ�
����*�3�a����3#����=�R}��<�]��_$��KJ5��-�zI�(��,&!�;������m5n����a�3��Q$�(QSg���&eu�{;�#mb6�=2��p?HZ��.J�R�
���ӫ-�Me����^�R�ʽR��U-�������$�'I;�IbN�wt�ĝ$��N)�t߂�HrAX�7�B�}���+�`����M�?7bP�B��o��[��<��s�aM���e_���'0lc��.�,k�}�a�/b���v'jI� 0,��{�|j�S�0�&��/�<j<J!�$��
�u6��믳lV�p��f>��u��Q&V�섪D��f���@8I$�Tk�hӳS^�k�h���]��B��w'fV\τ��8�ù�rI$��3����S�,w46�UR����;��nP����S����xxu��s��_H�\��W��6��CI$�eM��J�~�_SlQ���Z��'��ؽ"�z9�Ȯ����Hw�=�/�v�M����M�WEN���Y/Yb2dx ���14�g�-�2	��7�0��[�z��2T\�I'c'�{�}A����~܏)�T���t�B��L��fmp�FM��I$����C�Z�yr[�ZṊ��H>_�`˃0x��P�}p� ���/��<t����WX�f�3ͻ�Wί�σK��3������J�B�ҪQ�����+����QH�Qcb�0b"�"����
��J��D+l��D�$�PD%�K!����O���U�K.��U���/��r����{��%p�k�N:���5����te�m�z�2WbZ�ĖkP]�K�hJ-�
	��d@�1��I�Sq<�o/�n�q�t�f#�;�I-E$��$�����r/!z29��!��	 ������}�_���o VqY�zj(	1�fwD��ч�z6b܆|���͙�f`����Ǻ9�/z�r�����DK�q᣻1�ӄ�OZ��L=����ɓ�z��ԡW�>��b�Β�P�v�}����Wy�y�^�:}�CVI$�K��C�X�k��ҋ�S�T�E;�}�����#�H��~�����M>�I$�]�_K�.z�y���������_����r\�_�P��]�(~f`/�P'y_	)�9$���=��GC� H��|��=����6dE��zOQ���VZ~��#s�\we�����"�r�(I$������?Qʪd�ފ���+]��1�ֳ6e�1���G-�I$޷�+�.�q�)��x5Vκ����Wv�`qG�ո������!�$�ۺ�sƌQ�wƯ���VU�窄O�;�K�##x���HJ�g���QҶ#�Q$�aM��H�?i�WLҨ��Z�d�/���t���z$���iOy�"y{�I$�����Q��O�1��	�8�:�C��+]_[nN@5��tq�׃�4/q��ҳ.Q³��)����\�s�ްu��+1�$��4�@�_��G�:C�.��n��Mg3��gXڨo/H�y��v9�.S�h���ؗ�,��\��}����/��|�uWovq��$���wt�I����H$�蛌�v��m$�Y�G�d�d�K]��.��m�ZƤ��F��om�0fY�U�舕�J�r��mY$��n�6�t�x�E�X���\�LL�#7��w�	>}/��A!�$`����* R2{�0�
�m���Iw��v+0�:b�ס�^`����? �Rm��ɺ�	$�����a���t�1�����]��9*�j��������˔T¾�A��o;{2�s��ҷ�v�f
���3���.�-���Z������W����$��2��L غ��V_�9N����������υ>��D��˿A$�b����C����G�Suᒧ�S��5fx9_q�	��4N�{=�I$��2���[xa����E�Rx@w��}�����'UB�BI$�b�*(�J��WA����ĝz�/D/3=��i�ҕ�(˱�/3$�I�_8�з�f3�:24�õ<�Y�ٹ���r��c8����A`��UUTU��I
Y��BH`�x��p<P����p�>�s �H�`�UH���b�#ȁ �. �&RƔ\�院�M�!�Ny�Q������,0E"�" +��1`#"��dF*�B�DըȪ*�������Ub�#�te�*�RE(�7(�V��D�� �R�A� �A�A�5(,m��ƅ��A�bA*-oT?=:8���0�V�Yb[("bZ�03(6�Х�A2�h%�+A�J�,�4,��(�J4h6X��ZcYA���%�D�R�����A�JbŲ��R�Z�вб1�B�hR�,���д�iB��)B�V��ؔ���l�hZ"PD[Bʔ���e�bA�B��X�J62б�.nc��!eC��bD)JV��cYA��(ZX�Z( �,Tb$Q�PQD���E�ED�*ł1QX�"�"��`�,b"����Ŋ��PPX"DD`��,DX*�QQ�]�*�U�AA�,�b1U �1T�H�*#"�(����*"���?������H�E�(����PTF ���"*�Ȫ�E�`�Q`��PEEA***1F �����A�1c1dU�EQ ����Ag' ���A��Q�"��((e�0EA�PT�X��b�� **��UEV(��DH�1E��R��#���T�*UF1(�d�`�-eQTkFTPU�TE�
��X�9�O�h�E`2D 0Qb@Q��� 0PI! 
24�c$UP�X �U�D";��^,�A*&�DV)�����d�*��� 2z,�ђ�D��\3̸)������Vf��ݛtZ�eZ�3��4�L�1���,��@6Umd'���Z�e�g�_�I�<�o���C"��2���܊N�{O��������Ϩ��ý����8�bqӟ��S�����6��+!\��k�i�����?��`����Ǜa�<���p>�T$!�b8�[Lq�T�Ǽ��gSu�A{�.��=�*��wX�2ES?��1��:۽��ǘ��C�>�"P��4��Z=��n|��*���������\�����fc3x�7�"���Ƚ
�:�|�zC�@�#{��.XA���V�8���7���H|��g�D������eF��<�Uǵ�o=G������Z��T$���Liʼ"�(�0	�*ц�ʫC��&!��Ɋ�eLYK)b�U��'y����1�c%��1U�FYH�e��LĬ2�e&1V�b1�`MX} �̲(�f��1!�����F[�7:%8n��)T�n�B��AYaYPi  -��#>���fBk:s���B���W��E�j�ƶ��F��U�k����R�?��4�3m��]�įV����s{�L1D�d�)��OȤ���L����i؇�MɄRQ�Oq����Q����7o��������mn���s�_>1��c�<>[����M��q���9��]i�c���J��1h�mmc��Τ'ӂ�|����ä}����C�J]�<{�*�fk��U:-��xom#�>�"0�Qj�����ܪ��ߒyx��H��h:}rXu�"r"�I��XQ�3��~>�BNA�0�?Y���[� Cli���,-� ���
\ Si��X�Lj�J
���C�d���!w2*Q�2ȥ�J,��],371,����P��5 A�=~~Z�g���C��T�R��]'F����n�Ekl1�����g�ݴ=��}��ˬ>fE�B��*y�� ��H��R}A��y����$U:V��k�G�jf����܊�����J���������O�w�:{|��N�Q̆k�5���r�i1�W{�v�.\��O�7���/���!nhW�f��H��췿kus��;́��%�4ς���롘�8`m��
�I�		�4�ИM�b&��E2�I�<E���P�p�/s�ǁ�d��i�@ؑEQ�3m���f��7�wv�f'�Xmue�T��M��tμ}������\��b��<��qT��T�Z�q�i.mr��x�]$��6�T5�ߩN��o�C�*��2���．�yx[�U��H�
��� 