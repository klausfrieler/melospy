BZh91AY&SY�Ud� $w_�Py���g������`�}=�^�@ ���/���%T����@�  Z  � �@ ���(�
�4Sg�UT    �4�@ ��d��yG���� �Ʉh� �T��!F�hh�     zQL�d�      �B	��4�4��x�4�3D���DH�d¦ɔm4�)��  ���g1)��I"BtH!����$M@� �O���L�k�l�a$8� S,tk$�[m�ݴ�'\����ld�VI�&�x��~��f���K2"�,"�bɝ�ɡ������d",�h�IH�LҩD%R[l�C!F�F*$Q�Ui��
�C�USo͖ì��-�F�A+t��v�KO���,�F���T��I�\�(��JBJG�4M4�i����M�i�r�N<̐��*��4�l��IF�&�*�蜲���>m*�˪����;5V���Y�CR!4ij޷��flZ-t���P���6l[�E��S!�50���4h��Z�_�L�UБ"��С|���_"��:��(�y/��M�`�`e��g�3����P�8�9!W�oz�u��rVC�Ѯ��ȼ�;�\!!� $�N͖� �DС�fl�#�	�9�tu��y��"�o1�ŧۜ%�����a���Ж%&����h����4��G��2}"7{7#0Je͘�yM�͊k*�q]3d�#l�N����t���tnm	Z��Xܘ���i��Q&]H�ڠ��Nd\�>�37��vއ����{�o��Iٝ�8sj1=Z����܃)F勌�//sYM��N��
q�r�x%���h�os<��L\��)+�9[�H�*L�2�0��S �D1��iEahi�2H�-u��9%CAX(���$�Ɓ�Gb?�����|?m4�����������蝑��xx�,��w��-�;ţZ����*ZRa K��C8ILV��HZ-ln(�el̆Q��p��jME�C
�LI�^�TwsZ�D�ϱd��غ�nQ����p��i�Q�����J��$mҡ���FЃ��!\к�6or�����������7���@�u]#3j�����EP�O�@f�$�*5��]�)�OV��uh��m�E�[m�����ܜ�̩��X�7333v��$l؄�k	 	 !0��� ��S��!
@XL B` B�+��X��� �EQ'��vaТ�@D0�98{'�;)& 01���Ͻ~!�#$Oy��q�z��,_Nf��6�D�4(ͱ�ʔr�N�`Ԅ�B��e�/���b�P�RK\N���9��"uwv��A]yb�:�?Zx�akkI-��I$ǽ�g���j�D0���)��ڏN��"7u�q:��G��u{��S�FM)P��ɺ�B�,kb�tl����WēU/�ҊP����k\��L��rI�E#��LTN�q~Jsj��ت2"�
8�f�Y�y*���Uw����ȍ2d�&.dʹ�m:%����T�R2u�>�5Ͷ��MC~ŞՋ0�ᙀ�g�&#������bi�	��1�����7~��}8��?��N}�����m��m��PKX��fn��{G��k�Itqjb��HN���,�<���<�z1�Ç��M=��@�U�=�0z˪�#��:`��eD�Ӓdy��zio��zr�Z;y��[ DG�Y�M�G�D�*��-_Z��3�^i��Ny3kn�o�p^��4h��$pPЄ"&|�ځҦ���`P�2BI�ݏz�F�MpW�33�W��	��-�ҏ�k�A ���>H��ڢ0��ߩ��U>���@k���j1m����˖\fE�	b<D �|����fM(��nw��F�͈Ev��v��Ex0A'vF�)BQ����S�Ev�\�l.�t�p�t�6�U�S �G��#�9Ok��Պ/��/����w'�{�P6�P��X���d�c�p�ePn������u��s��;".������B��b�H@�ˆP��}b���9G�
c�}�b��="�uP��b ��G&/\�Π'c"04��1}:Fe�$B�nL�Ȱ%��ȉ�AȌFI�D�� ���׋�$�])@��fA�s�xq7 ���V]��W �%��ݞe�yts��z��̜=}ve��� �>$��Bsk:T�iU>s�`YGl�o����>��m��m��m�"^̱9�;���S=��^4�Û�j�f���5��UHLI! �[�w�q�4��ic���������z	���ic��W
��G��;c}��&fA�@,]C���f(=�1[:;#�*=$�� \p��Ԏ1���v�ӟ:�}�utN=�zm.$����S]��Ӻ�W��z�;�D�p�������oU��Ү��H��?�|��ać����#�_�ʛ�~��Y�7<q�F��Z���M*�j&�1����7���m��m��o�?��"=I�p���1߆�5����47�Iާ�$ҏS W�͹u@�H����4m�wNσ7Q�2�B��&}}@h�Ӥ�t��Vv���ԲH��+jh��8�T�"��@��  �G��z�Ze�@��D�-����`�^�^Ϭ��s7���*8��L�� ��lu��2���*��ׅ�5��U��:��$����G�ԅ(�3ED�,N�b�=[Q@罏�׳"	?!�$�zz2�z�bMJ☚�>��l�,����m��I$�2j�I=J�Yf"��b�!!I˸�V
��o������듺4����H`PHc���������;<�Ⱦb�j�}Y"h��P��F�@������n�+�w�1��:�}�]u�k�â�g:'�H�X!P�Dc�a\�\���[.E(�
�뭝�B�U;���R�8��v>�V�}A��/#P�2f{�ĕ��'Ï��Dx�}B�^v���ʋ�B�r�7&��b��n;�1dL٩+����E$dOQ��6�Y�wȍ^,���I$�I)b�� LzI�$�HgNY'�
�\zRSj�M�jy�D�`	��M3s��tPf�Ǉ�px�7=u��u��z� n��	�_Y��(G}c~���d�b1c g��3o%��輜@��4�<�긞^"QΑ8=1��߁1ۑ�t}������W���9sQt#�kV3������>�g�E�ؑs� �6�Q x�>��ٽ�K���^� �f�0-solH����&�r*[	*I$�I%�'���[W�١]��A��7o+�gi��,}�;��ܝ�#�څM>i�>��?V1Y���`�xD�$jo�L��l�еZ{>����N��\%�|(V��ӫ�`�1_)p������Q*lb������ݙ����Tn5����ӜЗ��6}	� L�=��ea�����/���
pP8D�yۺ����ىcQ��bx���@B�����H�I��`Mc)�J??W�	$�I$�I~Hb����?i���[Q��9t���D}Bjb�v_!�N�蠔i�RvEo�w�X٬��;g����2�9���3�3�w�w�2*���.
@��#��3��S�s�ol.;Y��[O�;Q�k�ZB�5Xb{M(F�32@p��J�< ��{�$p���cǞ��s^t'��b%Nl��M�uaX���rЦ9x��H${ď^��2&jk&�Y�qX��R�I$�IC���"��uw
���Q����3��-�m�X@D�D���W�*]�w��#�3�\C����GT�9Q�׳��! {�ۃ���K;So�\�G�<ؼ�{�<�����졘�O?qV�"A#)��&�e=Q/b����(T�ѥdI��Ma��x��a�28��
�~�u����=h���UU-�ڶ�m�TTD��SӤ8��@�coS*��Nd�8�Y'�(+�6�f�����
s�il�X��fI��)b��Z*�Uj�4Ѧ�V�e�Zh�,U*ʫ��jʶګ>��fѪ�4kT�K+��Uj֊2�K�D�9rL�v��\��X\YVL3%�V�afR�n�0��V�aqFe-\�:��Q��XVR��Q�IJŖ����Z,MX��Y0��&���6qb�d�bJY�aFU�%2d-ac,n�dh���Ն5��sF�i��t©�gM�*��L������R4f)LL�#,��I,�
f�jF�R�ZKD�ʡSy����f�mh�$ fBF)�Zh1RȪ�Y5"��Y�4|585�v2'���*{{l��)"IhH��"����r#�����e�e�oX�3L���
�wS5�+�A��ڣ��
g�6OH������Ȣ���#`��V����M��F�^n��?"K��N	��Px�f^T���A�8
����|�L��qn0y)�ӑ�� $�V1E|R���D[�"c�5���TP
�|��F�3ÚN��@A�r�tWh�
�r|ۗ���Dml��2���C���0��>y�3�9�9�"OK�w��z1ۼ
�P�I��C�-���
�T*��D��#�,�ie�,�[%UR-J�%��Y�-�*�T�!�X��ϴ&/=�9WIce!$E8�Vx%G0@}z�)�r���4IQ"�Ă�*���=$�����% ���*,�jbB�W`�h��u��hW�yA����=�1JIL��|����=����#���������,LN��f���m�d�U�� Z6h
�ң�&=�A�؜���t���[C�HI���X�1j`ι��=�	�l���V6O�Y #S���~A��� ��f�8I��T��W���/O�$�Sz\{�$�#%#�|���$8����,�=v�k���<�ɸD��"1��nD�q��Th����Yֶ�̪�"�d�G��+�Y�0���vJqQ��P���F8�����翮�8<�yE �Q[ހ��@h� ��3�t�;w�t�@��F��9�́���t(�Oq��\x戨@G�w�P1����?�f��QY��( �9��`D$5�	��tƊc��d��;���������]?^Po��e� 5�yF�up߆��P
�"����tv��1X��yNN�Rb�T�h��;�����'Y�X�=�&�0�ē����U#���<�
�����I� ��(iD@�ӷm��G!p
y��3�0<*E!z<��ewA�����A�뚇3
9y z0+��w$S�	�VL�