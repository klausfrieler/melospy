BZh91AY&SY���� Dw߀py����������`0�|��  �}�  r� �|����` �  �� 	4 ��` O@ �  �� 4    <�  O��4�JP����ک��� h   �   5<����M h     ��T
        M"�ҦQ�� ��   $�Si�z��OM'驓�M4 F��LL�QH&�Ѧ�����ʟ���e?Jh��h������D����oP�	"�@2.�?��߽� ^�*�
B�C�K��T����,@�*E�2� ��$�Q'G�d5�V�^��T�b#��da�LHD�!�#j}L:+�'���y�>�|=��r���}0$���X�(��m�Et�c�)�Y����:UYdL��suG�}D33�R4F�����b��d��ۨ���qv�5E2�e�b�ꢡiFL��nn��(�-�o`3fő���!�#\\�4p�f�����!��>e�p�D�Y���P�(� �D�-�w��B�����?5DQ��i=B�R�L��:���ZI�6�ȡIQC�JhY��!�2�cz�:B��C"H�L�r(�&�A��-ܕU[n����&�~DII�)�C2�{Z���Re�E���R�$A���X�HQ��Ɇ�U
"��T(��"��*��QE,�8�l:F��}$" �i��d�D�$L��?�Sv(�"ϙa����T(�d"�!N��P�� 2$0��d&��GZe��c8�ˎx��5556�.S)��o9�5
��8L�fgt�v���dnw�d�fÖ:�3im��T���w4�
E	u���E�9WK$&��AM*H|���N�j�6Nb
����)]ݣN��@�qC��N>��:Tcٜ�����sùq4cj�^��� �Dl�����$��G\��(ɽ0�I{���0/*���#I�9��'�+K�s	,�E��ō�~wt،���k&(ʧ0����,�U��/b�8�+*��
Z��$���Oh���3TD����u9�Q�M�j��Y6�f�-1�N;dt���kw˅�9�UN���i�F�a�����nJl�̉�*�)8�ΐ�P�8@A^O/I�� �B#oxH۸ш+Hp ̘�B�4��UDii�v1Ȫh#�+��L��`ۚ��2' ����*����;AlX2A�X�:攃N"��۴SJť�j �"�xh��hC��U���u�ԣ�-�ݬ�tn]D,t+0V��sQ�8�T�1Ef;��&Rn�a�%�:�e��ö��5pU2\6�����t�t����w:�C��*f/��"kra��.��TbM��n�$V,�^�ɚˈ��P��U�e�׶^+�qL���xY�x�%*@���'b�A�y�P�-��;{�ԻF���mPB*)����&C�5h�dn]dlļ�"����^;��n��[8��˺���ں�S3m�*j�ܻJ&�-n��G.�8m��-)r�U��h�e�L���)�����7n	��b�fֹG%�M���U�n涙2��ȕA5i)$�J
��eG�R
)���[�\̸UsZ�p�ͪ.4ʎ��㳏��:ӚGޞ�*���|*ح*�s��գQa���bs�erz��e'��̙�ś:�l���K���;�F�1��w��r�t�ֈja�S�"�0K��m0ݕ�$#LYb�# I���>���*Yle�+&�7q��FO�vkj��u.2��ݙv"e9h�v��Ӳ���.`Ū5[��1,Q�1�0g"��j�5��E�&-���92*�$T($M�t�ޜ��d���]ᨫ�3R']/7p��wb��r�����!�;�l�B���f��Nf�ʓ;nks-b,ВȨA��(Ld��P��t]Ί�����Q�QC*��ۻ���V�flU�J�(�&�FMg�~߸?�/���{��a�.W�hDm��Zi!$7���UUOMVn�uf�jjУ`�)k�Z� A�춽ً[;o��Ŧm3{a�{ݱ���k   `  A` 4�$�  $�U�F���T X 
  A  `  J�����VI#33,��A  ` � �\ 4� P@     ����;�;;����|nn<3�;+H#���N�t���Q���u/����/��*3�4km�1h�6�D��������uNQ��N
��GX��B�����/HZ���N�X�����x@#N\	 ɀ�]�L����Je7uj(f���kR�*���4K$[��Q�T̘%)�M�a�\��H,Qs]/�ܑx�]yj��k2\P�ݧ��zZ&M5J��BI$�3�BI$�;�;;�����ݤ���y�}�j�o(ǿc��d���|A .Oc�(�D�C�Te�Ы$����~�#k��鲲�-�nۭ�;j[&ۥX��6�qh�a�,V���k.�d�H�3u���RڡQ�j��D�ͣPW��a�95�g���fh��u�l�zE���"��՛���{�+j�zP5q����C��}QE�����ptdy�X�
�Ĕm���a��� A�"�ɦ*��$7&	b�r�$Xw�B���yN]ҒIBs"�y�T4C�p3`�}���55咠����I����,�؛VaΓ�̜��.��I:[r�"��S�c��{��'�"�X|C�"�VE;A��-m��T+E_	
�-�|������kJD~8�_����X�+��j3�6qӋ�WR������� |��S>���4ݬ" a��,�B!%�}a�U}����.��������{�X��^+�`�h�.Q�ȋN/�z� 9�>NW�C�#'cR��s#/XIHi�_�>����e��z�b���,C���xa�B�/s�e�j;(�ב`�}�3�����+�9+:d;�Ԥ���/6S��:F^�sh`������t�`��hM�6niS���ޒ�>�����=���:��ARV�2�t�(��E�q�G��{#)z�?@k��W3]T�c�_E8�jkyḐIj���ۍ͸jO4e����jo��j��x�7���{͌`�T����r�ս��rC~Ր嘃;P3�$��v�q-��+v@�H��e�(��ӫc1�F*V���~�:���5^}�sT<ĵih�*�NP��rg��DP6�h$+��ޛ({y� '�|EC��$T�2�8f�P����Z�����υB��&oi�J��T�Z��l���,���dY}U �	"��J\�cj56��/�����JP	L����7b#�:�l�6���Vt���۱wwwv.����#��I�R&�>E���&da�`��{�\�972n(����&C1�&�F[�K���L��7�k�ؚ��&N�Ogd�dI�ӹ#r�(�]��*�:�B�;u�B��۹�9o)�()ZlE��-�_kbh)&>������I�#V�2Y��U�8�0~1Vd�a��מ}T�`旼$������gM�
1��dG\z	>ص�6�t+ht!�o�:}�{�;c!}~w'6�)��A1���$ъE�>V��A��c��cLWqd������}��_b�l��KK�{�ZGѹ���a%�CWh_ �	���7���}7"f!�C?_����\��`ei*��zi-��?u@�)|
r��iB$�'����g	���"@�D�!��5V��V�7yx9�<�;�H8hrʱEdU��F���\��^{���H�'|� j�3����M�7��U��SX�j)���+sI���ƺ5�ȩƊ���\�4՛c�
�����)D$�I(������P��@��gT�|���C�-q�ݕ����5+U.���C,L1N�bP�p�N98�9�az�:��{�.W��#�ʡ��6s�(����&���d��6n�)�h�7���	H}��,�Pq��3�c8H�9{ã��u_������0���O�:��+��oLphmV`���%0�G��Q���MFl�u��7�2��0J�`Wt�_��:d� 7��WՈzH���ia�(,�C~?U�<�r9��p��Iq���Y �u���˔ZS'��a����fLWJ�̯*B�"��Tɯ��>��wV��!|b�)k;`p����rU꿎csծ8�94Dp��~^�SH����WF}�n�=���@�ގ�V{��1�P&.��tz_-��Ϫ7���Co>m��{l�j�[켰�\�uEϫ�	~��o��ղ`�ɪ�p!Zu�C([*�� �����Ê@��ƚh[��m��LۗH�;s�nE���S�W9bb�l�={+V3���&X����D���Ë3*��UY���L
�J2V!��bP�}�&�X=�c�os�P�&d��'l�%LU��4�Pa��'��xg��к��(�>����u'�t�R�C*�Ӡ>�id���׮r槢N\D�&�h۞�[,��Z�C��Q��R'"Ǻ���H��Ɵ1�^�8|#�GY:%�-X2:�����$5͒�ϼ�q���K���SZ���&u�^�S H|�S!��z�ʘ7��^�da9p�{?{�y��Cv�t ��gKn����������(i��U~��B#M�	$�q7����o�3�类,�mT���H�lA�| )��H���.朷�aR$�382'ޅ�&�)�z^�q}~I#���K��\/F�"B���> =�wb����=
)A��kq�A����G|υ��"�T��c�*"�("*��`��TPAQBj�r���5BI�%��7גvwJ����l��X���b���l�s�Ό��Ib��UT�gkڊαy}s�J9gS�逋���ay�1'G'������VWt;+�qb�����L��m�0�BHc5�X&6W����_2/����o���g�'�3�a�!VH�Bk���ۍ��ḳ�xP�p������5/hG������,�������*7�-g��=EgYn�kދ�X�5+�Hچn�ٻ����
���{fiH��)�H�
����5�Y�d@u���'���-|�iF����DzOW@��Ǉ� ���(��ޢ�V4F�u_Tijc�$ƭZwV{�ˍ��}3���&A>���ǩA0�G���\_�u�W�[.��O��2�I� F��b<���Dj�����#��N��y~��p��!�q�*Ɂ$�q"�[���͙�lD�R$���u+�j���(}5*�2�q�(��L�EY֌A>;���a��Q�-۫��l�-�ҩ��bc%�L�)%06[`�֑��0�ei�&��~����\S*���+�[;�k�̜�UU5��xxC�|�ʔ%	7j�RjR.t�T���٥���Z����?`�`�Cu��[�y�<>�[�+��.�ӧ=r����{�;b/����I�g�o������W�ӓ��&�7��Y@�R�w#�{����Oמ�N]ș� 7f1��1�F10�
�z�%k)�j���O�1���x^֌�Soܠ�^�$kx��w�� �	ɩ��2�����.k��x�bZ��lo��F����]�U�ʔ���j�������}���
�M:��> 	��9�|�헐����1�-�5O���NAK��=�<,���J��l���++��Z�	.�}S��w���^ݍ�E�9xxvvl�]�k��}��3���>'���'�h�����G�݅A�&\�Uj���b�rz}�H�X��AV(�PRG~�i�~��T��Li�F뷶�\�P�)C����T�^?!�II�-eq���ڢ���5^'���mͲvp��8I,%�9���3���)��� B�zz�dF���8�F:���}�^�#{c�hQK����B T���z:�w�P>$*G,��̎j'��y�~3�G��vo�'��1�W�_�>z�l��q����\��Ŭf'=u���ەr�2��!}�33&����?j�;���LXc9)צ�b�"xG�lw��mQ��p0L�>	T���������V�~P��������%Ck}\�n���{7/2�w\�E
P;�4]���;]�y��է3�*�m�D���];Yv�J�ȡ�֯���ơK�4�?�}?�8Vi�<3Ѩ� �,����"�랎u�k�<8��o"�#411n�l/����6M�V��qp^
.RH��/#	JS2d�IH3�PEJ2�3���(yIMd!&r�^d��y*��'�9M=��UU��]����د���������EI������'?�F�k�� g��iF�U�Ϸ��Kb�h�{�)�!sW�S��q�cڂ�Oܒ�sN����?�����џu}�}��y�u`��|��D.ڻ�� �3nc=�)�2Or���Ǥ�9@�·��s=b�s`���E�˱���D<�	�Y��q�_��}���i����g>NU����uJsc��E��wE��{���"s�}V�؎�{s֮�W������[u�j���Z5����J�gE���6��:r�>�Ȅx�)� 9Ȝ�"� �I�ׇܼj��Z��2'��	��*f{ǚ�b���PT��G�M�
2*��*��/��^E 	����av+Z�B*U�K��X�/Zt�"Q���!X4��ݮ�1s����ɣNEE`������WK#�_Mn֛����wwwV�1L-Z�^��U&�,�+ۋ�_%�5��l�Af�ț��'Q�~��/K�<K�pގ����}R������V6�T�i���'�	��'�� �C��k��=�6,B��T-�e���MA�GL��˪w!�������.�슎>ї{�7�c�lH�������3=�,�K��m˸��p:�x� �����#1w y\����97��,�F��c��	J��{�rM?����NYUf.�vwno\j/���D@�@
�qM�e@끗���%^f��c8��\A�d>�]1�/�@���,@�/��~����7��UT��Vť��ڶ��a���_v��3��)���>y�gL��à bd�M�
iƇF��3��3,�*id�����B�`�uh�cn+V[�(bb�d�21�(#�%��bœvO�X,i��cTs ���L1P���'��9�6#b��b(a,1��SQd���AU̗�#8d�`,Ra���9��
�"ᒀ-�1��@�#,d�(F�%BXʰdY,�΄*-�"��dP�,�
��2�����*�H62VE�ؒT��"
ì�a�!��"���$X,� X�PJ�E@V,�0������" �X��B((-�őHK**ARYJ�Y ��VIBأ `����!F,��$��%�f!D���!��P&L�*0	ch��
	Q �2D2��%����D��@�ؖH�Pj[�� (Yb4��lJ��xɣQ	cj�"���J4-��	u&L��)B�[�,��T@�-�b�#I�ٻs; d=�Y��
���bI�=��&����<�ZH�@�[!��2������m~�۸}�?}��:��D}�"լ��� I"�!�Om�S|g��� rG���?���NQ����'[ͯ�-�Ϳѡ$~j��b?���ԑ$pՐ����0+=�+,=�s#�C��Ľn	���Y�f=�V�S��lFh�R�>�W��3�i-��F��?i��	�"�%E*#ڍ$X�I�5��9�F��s��C�} �)1>���.������%PB�|�?=�oQ>\>�}��!	#!#-���$����tjþd���>��J��z3ͤN"�F�I#��NIa���oA�m�0G�����Z`��~"6f�(ˋv�S�cGT�q��=���=�'�%%�=m���~M;����W�dl�*h��	D�2�LSX�Y!e"�EE�QD�`�%��TP�Y$�,@ �H�6��IEB��*Ĳ�-�V%�AV%�ib&�Fx>�0]uaŋI��!A���Co1c��;�4'�QLY����( aT� �cd[
��;�\Z��spzS�~2Iia��qc�,����38�Gj�tn�$����$�'������#�k	�?M�f�c�ꊛbB$�m&I�͔���$�6��l�������$�bc�1��&Q=N3G�I�����j��%fi����сa�󪷛'�<���]���8z�_^��WH�$���Ql��[&;�J�?W�_��nɼ�6~���^ȎDW5H�s��ɶHI$Z�>�"I��4�O�|�N�C��\�e<X2�0��l��^pߺ�$�Rf�%����L����'�]�A�n���k�,����˯3��j�Γy��ޢ�"��I���!r`�8���I�Į3�%�,��J�a<ڐ��ܨa�x�g4��M#)2���:�3���mը�� H1QV��=�o�|B��:5;���T����7p(��Xk�j���/'��G�n~�5xu'͓.�ٗ�F�H�N�1\;x<eQ�Gqd�s��S�x��&�5��y����S�ׁ��G�䵕9N=��P�+I��0U!���C�o��{܎���x�;H�fφ�9����5�a�<����ѥi�`�b=���#9\�y�d�s��RJ�{u��3&�9�3S^����21��nl��A�""��ܺN�;P�oYe:vӤ�sY��5���������Rv8��,��n�7�dn��c�}CݩT��K:��"��j��g�ϴ��p�2������wϗ7˪u�i�"�k�
�`6�J��EMP�ȼ��<a����8���<����>���|E�$=͎�Xy�{����"�(Hl`�v�